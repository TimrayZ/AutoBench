module top_module (
	input [99:0] in,
	output reg [99:0] out
);


endmodule
