module top_module(
	input clk,
	input reset,
	input data,
	output start_shifting);


endmodule
