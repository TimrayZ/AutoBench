module top_module(
	input a, 
	input b,
	input c,
	output out
);


endmodule
