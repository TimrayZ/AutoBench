module top_module(
	input clk,
	input reset,
	output reg [9:0] q);


endmodule
