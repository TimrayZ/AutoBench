module top_module (
	input clk,
	input a, 
	output reg q
);


endmodule
