module top_module (
	input x3,
	input x2,
	input x1,
	output f
);


endmodule
