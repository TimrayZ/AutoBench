module top_module(
	input clk,
	input L,
	input q_in,
	input r_in,
	output reg Q);


endmodule
