module top_module (
	input d,
	input ena,
	output logic q
);


endmodule
