module top_module (
	input clk,
	input a, 
	output reg [2:0] q
);


endmodule
