module top_module (
	input a, 
	input b,
	input c,
	input d,
	output reg out
);


endmodule
