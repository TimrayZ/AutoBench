module top_module (
	input clk,
	input resetn,
	input x,
	input y,
	output f,
	output g
);


endmodule
