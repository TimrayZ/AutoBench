module top_module (
	input in,
	input [3:0] state,
	output reg [3:0] next_state,
	output out
);


endmodule
