module top_module(
	input [3:1] y,
	input w,
	output reg Y2);


endmodule
