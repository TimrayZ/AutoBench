module top_module (
	input clk,
	input reset,
	input x,
	output reg z
);


endmodule
