module top_module (
	input clk,
	input in,
	input reset,
	output [7:0] out_byte,
	output done
);


endmodule
