module top_module (
	input [3:0] in,
	output out_and,
	output out_or,
	output out_xor
);


endmodule
