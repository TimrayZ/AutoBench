module top_module(
	input clk, 
	input load, 
	input [9:0] data, 
	output tc
);


endmodule
