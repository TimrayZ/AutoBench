module top_module(
	input clk,
	input [7:0] in,
	output reg [7:0] pedge);


endmodule
