module top_module (
	input [5:0] y,
	input w,
	output Y1,
	output Y3
);


endmodule
