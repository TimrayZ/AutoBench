module top_module (
	input [7:0] in,
	output reg [2:0] pos
);


endmodule
