module top_module (
	input clk,
	input resetn,
	input in,
	output out
);


endmodule
