module top_module (
	input clk,
	input in,
	input reset,
	output done
);


endmodule
