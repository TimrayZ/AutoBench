module top_module(
	input ring, 
	input vibrate_mode,
	output ringer,
	output motor
);


endmodule
