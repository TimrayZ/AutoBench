module top_module(
	input clk,
	input reset,
	output [3:1] ena,
	output reg [15:0] q);


endmodule
