module top_module (
	input clk,
	input x,
	input [2:0] y,
	output reg Y0,
	output reg z
);


endmodule
