module top_module (
	input [254:0] in,
	output reg [7:0] out
);


endmodule
