module top_module (
	input a,
	input b,
	input c,
	input d,
	input e,
	output [24:0] out
);


endmodule
