module top_module (
	input [6:1] y,
	input w,
	output Y2,
	output Y4
);


endmodule
