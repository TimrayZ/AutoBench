module top_module (
	input [4:1] x,
	output logic f
);


endmodule
