module top_module (
	input clk,
	input in,
	input areset,
	output out
);


endmodule
