module top_module (
	input clk,
	input resetn,
	input [3:1] r,
	output [3:1] g
);


endmodule
