module top_module (
	input a,
	input b,
	input sel,
	output out
);


endmodule
