module top_module (
	input clk,
	input in,
	output logic out
);


endmodule
