module top_module(
	input clk,
	input load,
	input [255:0] data,
	output reg [255:0] q);


endmodule
