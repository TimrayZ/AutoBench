module top_module (
	input clk,
	input w,
	input R,
	input E,
	input L,
	output reg Q
);


endmodule
