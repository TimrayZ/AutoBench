module top_module (
	input clk,
	input j,
	input k,
	input reset,
	output out
);


endmodule
