module top_module(
	input clk,
	input reset,
	output shift_ena);


endmodule
