module top_module (
	input clk,
	input a,
	input b,
	output q,
	output state
);


endmodule
