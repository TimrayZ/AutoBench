module top_module (
	input clk,
	input reset,
	input in,
	output disc,
	output flag,
	output err);


endmodule
