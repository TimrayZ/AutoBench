module top_module (
	input clk,
	input j,
	input k,
	input areset,
	output out
);


endmodule
