module top_module (
	input clk,
	input d,
	input r,
	output logic q
);


endmodule
