module top_module (
	input [2:0] a, 
	output reg [15:0] q
);


endmodule
