module top_module (
	input clock,
	input a, 
	output reg p,
	output reg q
);


endmodule
