module top_module (
	input clk,
	input reset,
	input s,
	input w,
	output reg z
);


endmodule
