module top_module(
	input clk,
	input reset,
	output reg [3:0] q);


endmodule
