module top_module(
	input clk,
	input d,
	output reg q);


endmodule
