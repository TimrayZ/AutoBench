module top_module(
	input clk,
	input slowena,
	input reset,
	output reg [3:0] q);


endmodule
