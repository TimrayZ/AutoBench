module top_module(
	input clk,
	input reset,
	input [31:0] in,
	output reg [31:0] out);


endmodule
