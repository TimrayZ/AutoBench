module top_module(
	output one);


endmodule
