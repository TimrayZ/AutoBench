module top_module(
	input clk,
	input reset,
	output reg [31:0] q);


endmodule
