module top_module(
	input clk,
	input reset,
	output reg [4:0] q);


endmodule
