module top_module (
	input clk,
	input reset,
	input w,
	output z
);


endmodule
